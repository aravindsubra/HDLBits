module top_module ( input a, input b, output out );
    mod_a u(a, b, out);
endmodule
